// `include "spc700.vh"

import spc700::*;

module SPC700_MCode(
    input CLK,
    input RST_N,
    input EN,
    input [7:0] IR,
    input [3:0] STATE,
    output MCode_r M
);

// 31 bits
//   stateCtrl,  addrCtrl, regMode, regAXY,        ALUCtrl,  outBus
//         addrBus                        busCtrl
localparam MicroInst_r M_TAB[0:4095] = '{
	// 00 NOP
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 01 TCALL 0
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101},// ['PCH->[SP]', 'SP//']
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100},// ['PCL->[SP]', 'SP//']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]->DR']
	{2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]:DR->PC']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 02 SET1 d.0
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010110,3'b000},// ['ALU{[AX]|01}', 'ALU{}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 03 BBS d.0
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 04 OR A, d
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000100,3'b000},// ['ALU{A|[AX]}', 'ALU{}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 05 OR A, !a
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'PC++']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000100,3'b000},// ['ALU{A|[AX]}', 'ALU{}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},	
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 06 OR A, {X}
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100101,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['X->AL', 'P->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000100,3'b000},// ['ALU{A|[AX]}', 'ALU{}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 07 OR A, {d+X}
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+X->AL']
	{2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR', 'AL+1->AL']
	{2'b00,2'b01,6'b011010,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->AH', 'DR->AL']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000100,3'b000},// ['ALU{A|[AX]}', 'ALU{}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 08 OR #i
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00010,2'b01,5'b00000,6'b000100,3'b000},// ['ALU{A|[PC]}', 'ALU{}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 09 OR dd, ds
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00110,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->T']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b01100,6'b000100,3'b000},// ['ALU{T|[AX]}', 'ALU{}->T', 'Flags']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 0A OR1 C, m.b
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]&1F->AH', '[PC]->DR', 'PC++']
	{2'b10,2'b01,6'b000000,5'b01010,2'b00,5'b10111,6'b011001,3'b000},// ['ALU{C|[AX].b}', 'ALU{}->C']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 0B ASL d
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b00000,6'b001010,3'b000},// ['ALU{[AX]<<1}', 'ALU{}->T', 'Flags']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 0C ASL !a
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b00000,6'b001010,3'b000},// ['ALU{[AX]<<1}', 'ALU{}->T', 'Flags']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},	
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 0D PUSH PSW
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b10,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b011},// ['PSW->[SP]']
	{2'b10,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b000},// ['SP//']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 0E TSET1 !a
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00011,2'b00,5'b00000,6'b000101,3'b000},// ['ALU{[AX]}', 'Flags']
	{2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b00000,6'b001111,3'b000},// ['ALU{[AX]|A}', 'ALU{}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 0F BRK
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b01111,2'b00,5'b00000,6'b000000,3'b000},// ['1->B']
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101},// ['PCH->[SP]', 'SP//']
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100},// ['PCL->[SP]', 'SP//']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b011},// ['PSW->[SP]', 'SP//']
	{2'b00,2'b00,6'b000000,5'b01000,2'b00,5'b00000,6'b000000,3'b000},// ['0->I']
	{2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]->DR']
	{2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]:DR->PC']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 10 BPL
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR, 'PC++'']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 11 TCALL 1
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101},// ['PCH->[SP]', 'SP//']
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100},// ['PCL->[SP]', 'SP//']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]->DR']
	{2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]:DR->PC']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 12 CLR1 d.0
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010101,3'b000},// ['ALU{[AX]&~01}', 'ALU{}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 13 BBC d.0
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 14 OR A, d+X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+X->AL']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000100,3'b000},// ['ALU{A|[AX]}', 'ALU{}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 15 OR A, !a+X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b011000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'AL+X->AL', 'PC++']
	{2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AH+Carry->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000100,3'b000},// ['ALU{A|[AX]}', 'ALU{}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 16 OR A, !a+Y
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b011001,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'AL+Y->AL', 'PC++']
	{2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AH+Carry->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000100,3'b000},// ['ALU{A|[AX]}', 'ALU{}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},	
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 17 OR A, {d}+Y
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR', 'AL+1->AL']
	{2'b00,2'b01,6'b011011,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->AH', 'DR+Y->AL']
	{2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AH+Carry->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000100,3'b000},// ['ALU{A|[AX]}', 'ALU{}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 18 OR d, #i
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00101,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->T', 'PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000100,3'b000},// ['ALU{T|[AX]}', 'ALU{}->T', 'Flags']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 19 OR {X}, {Y}
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100110,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['Y->AL', 'P->AH']
	{2'b00,2'b01,6'b100101,5'b00110,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->T', 'X->AL', 'P->AH']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000100,3'b000},// ['ALU{T|[AX]}', 'ALU{}->T', 'Flags']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 1A DECW d
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000010,3'b000},// ['ALU{[AX]-1}', 'ALU{}->T']
	{2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]', 'AL+1->AL']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000001,3'b000},// ['ALU{[AX]-C}', 'ALU{}->T', 'Flags']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},	
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 1B ASL d+X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+X->AL']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b00000,6'b001010,3'b000},// ['ALU{[AX]<<1}', 'ALU{}->T', 'Flags']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 1C ASL A
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00011,2'b01,5'b00001,6'b001010,3'b000},// ['ALU{A<<1}', 'ALU{}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 1D DEC X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00011,2'b10,5'b00101,6'b000010,3'b000},// ['ALU{X-1}', 'ALU{}->X', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 1E CMP X, !a
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'PC++']
	{2'b10,2'b01,6'b000000,5'b00011,2'b00,5'b00100,6'b010011,3'b000},// ['ALU{X-[AX]}', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 1F JMP [!a+X]
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b011000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'AL+X->AL', 'PC++']
	{2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AH+Carry->AH']
	{2'b00,2'b01,6'b111100,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR', 'AX+1->AX']
	{2'b10,2'b01,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]:DR->PC']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 20 CLRP
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b01000,2'b00,5'b00000,6'b000000,3'b000},// ['Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 21 TCALL 2
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101},// ['PCH->[SP]', 'SP//']
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100},// ['PCL->[SP]', 'SP//']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]->DR']
	{2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]:DR->PC']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 22 SET1 d.1
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010110,3'b000},// ['ALU{[AX]|02}', 'ALU{}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 23 BBS d.1
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 24 AND A, d
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000101,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 25 AND A, !a
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'PC++']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000101,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 26 AND A, {X}
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100101,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['X->AL', 'P->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000101,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 27 AND A, {d+X}
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+X->AL']
	{2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR', 'AL+1->AL']
	{2'b00,2'b01,6'b011010,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->AH', 'DR->AL']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000101,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 28 AND #i
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00010,2'b01,5'b00000,6'b000101,3'b000},// ['ALU{[PC]}->A', 'PC++', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 29 AND dd, ds
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00110,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->T']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000101,3'b000},// ['ALU{[AX]}->T', 'Flags']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 2A OR1 C, !m.b
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'PC++']
	{2'b10,2'b01,6'b000000,5'b01010,2'b00,5'b10111,6'b011001,3'b000},// ['ALU{C|~[AX].b}', 'ALU{}->C']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},	
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 2B ROL d
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b00000,6'b001100,3'b000},// ['ALU{[AX]}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 2C ROL !a
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b001100,3'b000},// ['ALU{[AX]}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 2D PUSH A
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b10,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b001},// ['A->[SP]']
	{2'b10,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b000},// ['SP//']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 2E CBNE d, r
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b010011,3'b000},// ['ALU{[AX]}']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 2F BRA
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 30 BMI
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 31 TCALL 3
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101},// ['PCH->[SP]', 'SP//']
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100},// ['PCL->[SP]', 'SP//']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]->DR']
	{2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]:DR->PC']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 32 CLR1 d.1
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010101,3'b000},// ['ALU{[AX]&~02}', 'ALU{}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 33 BBC d.1
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 34 AND A, d+X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+X->AL']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000101,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 35 AND A, !a+X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b011000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'AL+X->AL', 'PC++']
	{2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AH+Carry->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000101,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 36 AND A, !a+Y
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b011001,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'AL+Y->AL', 'PC++']
	{2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AH+Carry->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000101,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},	
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 37 AND A, {d}+Y
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR', 'AL+1->AL']
	{2'b00,2'b01,6'b011011,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->AH', 'DR+Y->AL']
	{2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AH+Carry->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000101,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 38 AND d, #i
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00101,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->T', 'PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000101,3'b000},// ['ALU{[AX]}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 39 AND {X}, {Y}
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100110,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['Y->AL', 'P->AH']
	{2'b00,2'b01,6'b100101,5'b00110,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->T', 'X->AL', 'P->AH']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000101,3'b000},// ['ALU{[AX]}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 3A INCW d
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000011,3'b000},// ['ALU{[AX]+1}', 'ALU{}->T']
	{2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]', 'AL+1->AL']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b001001,3'b000},// ['ALU{[AX]+C}', 'ALU{}->T', 'Flags']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 3B ROL d+X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+X->AL']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b00000,6'b001100,3'b000},// ['ALU{[AX]}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},	
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 3C ROL A
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00011,2'b01,5'b00001,6'b001100,3'b000},// ['ALU{A}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 3D INC X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00011,2'b10,5'b00101,6'b000011,3'b000},// ['ALU{X}->X', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 3E CMP X, d
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b10,2'b01,6'b000000,5'b00011,2'b00,5'b00100,6'b010011,3'b000},// ['ALU{X-[AX]}', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 3F CALL !a
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'PC++']
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101},// ['PCH->[SP]', 'SP//']
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100},// ['PCL->[SP]', 'SP//']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b10,2'b00,6'b000000,5'b01110,2'b00,5'b00000,6'b000000,3'b000},// ['AX->PC']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 40 SETP
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b01000,2'b00,5'b00000,6'b000000,3'b000},// ['Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 41 TCALL 4
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101},// ['PCH->[SP]', 'SP//']
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100},// ['PCL->[SP]', 'SP//']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]->DR']
	{2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]:DR->PC']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 42 SET1 d.2
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010110,3'b000},// ['ALU{[AX]|04}', 'ALU{}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 43 BBS d.2
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 44 EOR A, d
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000110,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 45 EOR A, !a
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'PC++']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000110,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 46 EOR A, {X}
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100101,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['X->AL', 'P->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000110,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 47 EOR A, {d+X}
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+X->AL']
	{2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR', 'AL+1->AL']
	{2'b00,2'b01,6'b011010,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->AH', 'DR->AL']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000110,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 48 EOR #i
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00010,2'b01,5'b00000,6'b000110,3'b000},// ['ALU{[PC]}->A', 'PC++', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 49 EOR dd, ds
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00110,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->T']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000110,3'b000},// ['ALU{[AX]}->T', 'Flags']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 4A AND1 C, m.b
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]&1F->AH', '[PC]->DR', 'PC++']
	{2'b10,2'b01,6'b000000,5'b01010,2'b00,5'b10111,6'b010111,3'b000},// ['ALU{[AX]}->C']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 4B LSR d
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b00000,6'b001011,3'b000},// ['ALU{[AX]}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 4C LSR !a
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b001011,3'b000},// ['ALU{[AX]}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 4D PUSH X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b10,6'b000000,5'b00000,2'b00,5'b00100,6'b000000,3'b001},// ['X->[SP]']
	{2'b10,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b000},// ['SP//']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 4E TCLR1 !a
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00011,2'b00,5'b00000,6'b000101,3'b000},// ['ALU{[AX]}', 'Flags']
	{2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b00000,6'b001110,3'b000},// ['ALU{[AX]}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 4F PCALL u
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101},// ['PCH->[SP]', 'SP//']
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100},// ['PCL->[SP]', 'SP//']
	{2'b10,2'b00,6'b000000,5'b10010,2'b00,5'b00000,6'b000000,3'b000},// ['FF:AL->PC']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 50 BVC
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 51 TCALL 5
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101},// ['PCH->[SP]', 'SP//']
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100},// ['PCL->[SP]', 'SP//']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]->DR']
	{2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]:DR->PC']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 52 CLR1 d.2
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010101,3'b000},// ['ALU{[AX]&~04}', 'ALU{}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 53 BBC d.2
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 54 EOR A, d+X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+X->AL']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000110,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 55 EOR A, !a+X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b011000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'AL+X->AL', 'PC++']
	{2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AH+Carry->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000110,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 56 EOR A, !a+Y
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b011001,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'AL+X->AL', 'PC++']
	{2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AH+Carry->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000110,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},	
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 57 EOR A, {d}+Y
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR', 'AL+1->AL']
	{2'b00,2'b01,6'b011011,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->AH', 'DR+Y->AL']
	{2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AH+Carry->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000110,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 58 EOR d, #i
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00101,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->T', 'PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000110,3'b000},// ['ALU{[AX]}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 59 EOR {X}, {Y}
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100110,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['Y->AL', 'P->AH']
	{2'b00,2'b01,6'b100101,5'b00110,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->T', 'X->AL', 'P->AH']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000110,3'b000},// ['ALU{[AX]}->T', 'Flags']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 5A CMPW YA, d
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00011,2'b00,5'b00000,6'b010011,3'b000},// ['ALU{A-[AX]}']
	{2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+1->AL']
	{2'b10,2'b01,6'b000000,5'b00011,2'b00,5'b01000,6'b010000,3'b000},// ['ALU{[AX]}', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 5B LSR d+X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+X->AL']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b00000,6'b001011,3'b000},// ['ALU{[AX]}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 5C LSR A
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00011,2'b01,5'b00001,6'b001011,3'b000},// ['ALU{A}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 5D MOV X, A
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00011,2'b10,5'b00001,6'b000000,3'b000},// ['ALU{A}->X', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 5E CMP Y, !a
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'PC++']
	{2'b10,2'b01,6'b000000,5'b00011,2'b00,5'b01000,6'b010011,3'b000},// ['ALU{Y-[AX]}', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 5F JMP !a
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b10,2'b00,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]:DR->PC']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 60 CLRC
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b01000,2'b00,5'b00000,6'b000000,3'b000},// ['Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 61 TCALL 6
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101},// ['PCH->[SP]', 'SP//']
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100},// ['PCL->[SP]', 'SP//']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]->DR']
	{2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]:DR->PC']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 62 SET1 d.3
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010110,3'b000},// ['ALU{[AX]|08}', 'ALU{}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 63 BBS d.3
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 64 CMP A, d
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b10,2'b01,6'b000000,5'b00011,2'b00,5'b00000,6'b010011,3'b000},// ['ALU{A-[AX]}', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 65 CMP A, !a
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'PC++']
	{2'b10,2'b01,6'b000000,5'b00011,2'b00,5'b00000,6'b010011,3'b000},// ['ALU{A-[AX]}', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 66 CMP A, {X}
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100101,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['X->AL', 'P->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b00,5'b00000,6'b010011,3'b000},// ['ALU{A-[AX]}', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 67 CMP A, {d+X}
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+X->AL']
	{2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR', 'AL+1->AL']
	{2'b00,2'b01,6'b011010,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->AH', 'DR->AL']
	{2'b10,2'b01,6'b000000,5'b00011,2'b00,5'b00000,6'b010011,3'b000},// ['ALU{A-[AX]}', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 68 CMP #i
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00010,2'b00,5'b00000,6'b010011,3'b000},// ['ALU{A-[PC]}', 'PC++', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 69 CMP dd, ds
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00110,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->T']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b010011,3'b000},// ['ALU{[AX]-T}', 'Flags']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// 
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 6A AND1 C, !m.b
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', '[PC]->DR', 'PC++']
	{2'b10,2'b01,6'b000000,5'b01010,2'b00,5'b10111,6'b011000,3'b000},// ['ALU{[AX]}->C']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 6B ROR d
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b00000,6'b001101,3'b000},// ['ALU{[AX]}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 6C ROR !a
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b001101,3'b000},// ['ALU{[AX]}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 6D PUSH Y
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b10,6'b000000,5'b00000,2'b00,5'b01000,6'b000000,3'b001},// ['Y->[SP]']
	{2'b10,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b000},// ['SP//']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 6E DBNZ d, r
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000010,3'b000},// ['ALU{[AX]}->T']
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b01101,6'b000000,3'b001},// ['T->[AX]']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 6F RET
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b10000,2'b00,5'b00000,6'b000000,3'b000},// ['SP++']
	{2'b00,2'b10,6'b000000,5'b10000,2'b00,5'b00000,6'b000000,3'b000},// ['[SP]->DR', 'SP++']
	{2'b00,2'b10,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000},// ['[SP]:DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 70 BVS
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 71 TCALL 7
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101},// ['PCH->[SP]', 'SP//']
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100},// ['PCL->[SP]', 'SP//']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]->DR']
	{2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]:DR->PC']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 72 CLR1 d.3
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010101,3'b000},// ['ALU{[AX]&~08}', 'ALU{}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 73 BBC d.3
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 74 CMP A, d+X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+X->AL']
	{2'b10,2'b01,6'b000000,5'b00011,2'b00,5'b00000,6'b010011,3'b000},// ['ALU{A-[AX]}', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 75 CMP A, !a+X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b011000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'AL+X->AL', 'PC++']
	{2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AH+Carry->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b00,5'b00000,6'b010011,3'b000},// ['ALU{A-[AX]}', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 76 CMP A, !a+Y
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b011001,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'AL+X->AL', 'PC++']
	{2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AH+Carry->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b00,5'b00000,6'b010011,3'b000},// ['ALU{A-[AX]}', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 77 CMP A, {d}+Y
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR', 'AL+1->AL']
	{2'b00,2'b01,6'b011011,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->AH', 'DR+Y->AL']
	{2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AH+Carry->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b00,5'b00000,6'b010011,3'b000},// ['ALU{A-[AX]}', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 78 CMP d, #i
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00101,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->T', 'PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b010011,3'b000},// ['ALU{[AX]-T}', 'Flags']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// 
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 79 CMP {X}, {Y}
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100110,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['Y->AL', 'P->AH']
	{2'b00,2'b01,6'b100101,5'b00110,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->T', 'X->AL', 'P->AH']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b010011,3'b000},// ['ALU{[AX]-T}', 'Flags']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// 
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 7A ADDW YA, d
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b010001,3'b000},// ['ALU{[AX]}->A']
	{2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+1->AL']
	{2'b10,2'b01,6'b000000,5'b00011,2'b11,5'b01000,6'b010010,3'b000},// ['ALU{[AX]}->Y']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 7B ROR d+X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+X->AL']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b00000,6'b001101,3'b000},// ['ALU{[AX]}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 7C ROR A
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00011,2'b01,5'b00001,6'b001101,3'b000},// ['ALU{A}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 7D MOV A, X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00011,2'b01,5'b00101,6'b000000,3'b000},// ['ALU{X}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 7E CMP Y, d
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b10,2'b01,6'b000000,5'b00011,2'b00,5'b01000,6'b010011,3'b000},// ['ALU{Y-[AX]}', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 7F RETI
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b10000,2'b00,5'b00000,6'b000000,3'b000},// ['SP++']
	{2'b00,2'b10,6'b000000,5'b10001,2'b00,5'b00000,6'b000000,3'b000},// ['[SP]->PSW']
	{2'b00,2'b00,6'b000000,5'b10000,2'b00,5'b00000,6'b000000,3'b000},// ['SP++']
	{2'b00,2'b10,6'b000000,5'b10000,2'b00,5'b00000,6'b000000,3'b000},// ['[SP]->DR', 'SP++']
	{2'b10,2'b10,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000},// ['[SP]:DR->PC']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 80 SETC
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b01000,2'b00,5'b00000,6'b000000,3'b000},// ['Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 81 TCALL 8
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101},// ['PCH->[SP]', 'SP//']
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100},// ['PCL->[SP]', 'SP//']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]->DR']
	{2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]:DR->PC']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 82 SET1 d.4
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010110,3'b000},// ['ALU{[AX]|10}', 'ALU{}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 83 BBS d.4
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 84 ADC A, d
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000111,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 85 ADC A, !a
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'PC++']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000111,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 86 ADC A, {X}
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100101,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['X->AL', 'P->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000111,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 87 ADC A, {d+X}
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+X->AL']
	{2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR', 'AL+1->AL']
	{2'b00,2'b01,6'b011010,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->AH', 'DR->AL']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000111,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 88 ADC #i
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00010,2'b01,5'b00000,6'b000111,3'b000},// ['ALU{[PC]}->A', 'PC++', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 89 ADC dd, ds
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00110,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->T']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000111,3'b000},// ['ALU{[AX]}->T', 'Flags']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 8A EOR1 C, m.b
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]&1F->AH', '[PC]->DR', 'PC++']
	{2'b10,2'b01,6'b000000,5'b01010,2'b00,5'b10111,6'b011011,3'b000},// ['ALU{[AX]}->C']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 8B DEC d
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000010,3'b000},// ['ALU{[AX]-1}', 'ALU{}->T', 'Flags']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 8C DEC !a
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000010,3'b000},// ['ALU{[AX]-1}', 'ALU{}->T', 'Flags']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 8D MOV Y, #i
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00010,2'b11,5'b00000,6'b000000,3'b000},// ['ALU{[PC]}->Y', 'PC++', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 8E POP PSW
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b10000,2'b00,5'b00000,6'b000000,3'b000},// ['SP++']
	{2'b00,2'b10,6'b000000,5'b10001,2'b00,5'b00000,6'b000000,3'b000},// ['[SP]->PSW']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 8F MOV d, #i
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00101,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->T', 'PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 90 BCC
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 91 TCALL 9
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101},// ['PCH->[SP]', 'SP//']
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100},// ['PCL->[SP]', 'SP//']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]->DR']
	{2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]:DR->PC']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 92 CLR1 d.4
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010101,3'b000},// ['ALU{[AX]&~10}', 'ALU{}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 93 BBC d.4
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 94 ADC A, d+X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+X->AL']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000111,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 95 ADC A, !a+X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b011000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'AL+X->AL', 'PC++']
	{2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AH+Carry->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000111,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 96 ADC A, !a+Y
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b011001,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'AL+X->AL', 'PC++']
	{2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AH+Carry->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000111,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 97 ADC A, {d}+Y
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR', 'AL+1->AL']
	{2'b00,2'b01,6'b011011,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->AH', 'DR+Y->AL']
	{2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AH+Carry->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000111,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 98 ADC d, #i
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00101,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->T', 'PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000111,3'b000},// ['ALU{[AX]}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 99 ADC {X}, {Y}
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100110,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['Y->AL', 'P->AH']
	{2'b00,2'b01,6'b100101,5'b00110,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->T', 'X->AL', 'P->AH']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000111,3'b000},// ['ALU{[AX]}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 9A SUBW YA, d
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b010011,3'b000},// ['ALU{[AX]}->A']
	{2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+1->AL']
	{2'b10,2'b01,6'b000000,5'b00011,2'b11,5'b01000,6'b010100,3'b000},// ['ALU{[AX]}->Y']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 9B DEC d+X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+X->AL']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000010,3'b000},// ['ALU{[AX]-1}', 'ALU{}->T', 'Flags']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 9C DEC A
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00011,2'b01,5'b00001,6'b000010,3'b000},// ['ALU{A-1}', 'ALU{}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 9D MOV X, SP
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00011,2'b10,5'b11101,6'b000000,3'b000},// ['ALU{SP}->X', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 9E DIV YA, X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100001,3'b000},// ['ALU{YA/X}']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100001,3'b000},// ['ALU{YA/X}']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100001,3'b000},// ['ALU{YA/X}']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100001,3'b000},// ['ALU{YA/X}']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100001,3'b000},// ['ALU{YA/X}']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100001,3'b000},// ['ALU{YA/X}']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100001,3'b000},// ['ALU{YA/X}']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100001,3'b000},// ['ALU{YA/X}']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100001,3'b000},// ['ALU{YA/X}']
	{2'b00,2'b00,6'b000000,5'b00011,2'b01,5'b11001,6'b100001,3'b000},// ['ALU{YA/X}']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['ALU{}->YA', 'ALU{YA/X}', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// 9F XCN
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00011,2'b01,5'b00001,6'b011101,3'b000},// ['ALU{A}->A', 'Flags']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},	
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	//A0 EI
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b01000,2'b00,5'b00000,6'b000000,3'b000},// ['Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// A1 TCALL 10
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101},// ['PCH->[SP]', 'SP//']
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100},// ['PCL->[SP]', 'SP//']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]->DR']
	{2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]:DR->PC']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// A2 SET1 d.5
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010110,3'b000},// ['ALU{[AX]|20}', 'ALU{}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// A3 BBS d.5
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// A4 SBC A, d
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b001000,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// A5 SBC A, !a
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'PC++']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b001000,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// A6 SBC A, {X}
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100101,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['X->AL', 'P->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b001000,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// A7 SBC A, {d+X}
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+X->AL']
	{2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR', 'AL+1->AL']
	{2'b00,2'b01,6'b011010,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->AH', 'DR->AL']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b001000,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// A8 SBC #i
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00010,2'b01,5'b00000,6'b001000,3'b000},// ['ALU{[PC]}->A', 'PC++', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// A9 SBC dd, ds
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00110,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->T']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b001000,3'b000},// ['ALU{[AX]}->T', 'Flags']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// AA MOV1 C, m.b
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]&1F->AH', '[PC]->DR', 'PC++']
	{2'b10,2'b01,6'b000000,5'b01010,2'b00,5'b00011,6'b000000,3'b000},// ['ALU{[AX]}->C']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// AB INC d
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000011,3'b000},// ['ALU{[AX]}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// AC INC !a
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000011,3'b000},// ['ALU{[AX]}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// AD CMP Y, #i
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00010,2'b00,5'b01000,6'b010011,3'b000},// ['ALU{Y-[PC]}, 'PC++', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},	
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// AE POP A
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b10000,2'b00,5'b00000,6'b000000,3'b000},// ['SP++']
	{2'b00,2'b10,6'b000000,5'b00000,2'b01,5'b00000,6'b000000,3'b000},// ['[SP]->A']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// AF MOV {X}+, A
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100101,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['X->AL', 'P->AH']
	{2'b00,2'b00,6'b000000,5'b00000,2'b10,5'b00101,6'b000011,3'b000},// ['X++']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b001},// ['A->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// B0 BCS
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// B1 TCALL 11
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101},// ['PCH->[SP]', 'SP//']
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100},// ['PCL->[SP]', 'SP//']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]->DR']
	{2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]:DR->PC']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// B2 CLR1 d.5
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010101,3'b000},// ['ALU{[AX]&~20}', 'ALU{}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// B3 BBC d.5
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// B4 SBC A, d+X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+X->AL']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b001000,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// B5 SBC A, !a+X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b011000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'AL+X->AL', 'PC++']
	{2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AH+Carry->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b001000,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// B6 SBC A, !a+Y
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b011001,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'AL+X->AL', 'PC++']
	{2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AH+Carry->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b001000,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// B7 SBC A, {d}+Y
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR', 'AL+1->AL']
	{2'b00,2'b01,6'b011011,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->AH', 'DR+Y->AL']
	{2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AH+Carry->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b001000,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// B8 SBC d, #i
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00101,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->T', 'PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b001000,3'b000},// ['ALU{[AX]}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// B9 SBC {X}, {Y}
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100110,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['Y->AL', 'P->AH']
	{2'b00,2'b01,6'b100101,5'b00110,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->T', 'X->AL', 'P->AH']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b001000,3'b000},// ['ALU{[AX]}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// BA MOV YA, d
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000000,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'b00,2'b00,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+1->AL']
	{2'b10,2'b01,6'b000000,5'b00011,2'b11,5'b00000,6'b000000,3'b000},// ['ALU{[AX]}->Y', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// BB INC d+X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+X->AL']
	{2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000011,3'b000},// ['ALU{[AX]}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// BC INC A
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00011,2'b01,5'b00001,6'b000011,3'b000},// ['ALU{A}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// BD MOV SP, X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00100,2'b00,5'b00000,6'b000000,3'b000},// ['X->SP']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// BE DAS
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00111,2'b01,5'b00000,6'b011111,3'b000},// ['ALU{A}->A', 'Flags']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// BF MOV A, {X}+
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100101,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['X->AL', 'P->AH']
	{2'b00,2'b00,6'b000000,5'b00000,2'b10,5'b00101,6'b000011,3'b000},// ['X++']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000000,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// C0 DI
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b01000,2'b00,5'b00000,6'b000000,3'b000},// ['Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},	
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// C1 TCALL 12
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101},// ['PCH->[SP]', 'SP//']
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100},// ['PCL->[SP]', 'SP//']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]->DR']
	{2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]:DR->PC']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// C2 SET1 d.6
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010110,3'b000},// ['ALU{[AX]|40}', 'ALU{}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// C3 BBS d.6
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// C4 MOV d, A
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b001},// ['A->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// C5 MOV !a, A
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b001},// ['A->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// C6 MOV {X}, A
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100101,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['X->AL', 'P->AH']
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b001},// ['A->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// C7 MOV {d+X}, A
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+X->AL']
	{2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR', 'AL+1->AL']
	{2'b00,2'b01,6'b011010,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->AH', 'DR->AL']
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b001},// ['A->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// C8 CMP X, #i
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00010,2'b00,5'b00100,6'b010011,3'b000},// ['ALU{X-[PC]}', 'PC++', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},	
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// C9 MOV !a, X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00100,6'b000000,3'b001},// ['X->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// CA MOV1 m.b, C
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]&1F->AH', '[PC]->DR', 'PC++']
	{2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010101,3'b000},// ['ALU{[AX]}->T']
	{2'b00,2'b00,6'b000000,5'b01011,2'b00,5'b11111,6'b010110,3'b000},// ['ALU{T}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// CB MOV d, Y
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01000,6'b000000,3'b001},// ['Y->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// CC MOV !a, Y
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01000,6'b000000,3'b001},// ['Y->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// CD MOV X, #i
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00010,2'b10,5'b00000,6'b000000,3'b000},// ['ALU{[PC]}->X', 'PC++', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// CE POP X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b10000,2'b00,5'b00000,6'b000000,3'b000},// ['SP++']
	{2'b00,2'b10,6'b000000,5'b00000,2'b10,5'b00000,6'b000000,3'b000},// ['[SP]->X']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// CF MUL YA
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100000,3'b000},// ['ALU{Y*A}']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100000,3'b000},// ['ALU{Y*A}']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100000,3'b000},// ['ALU{Y*A}']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100000,3'b000},// ['ALU{Y*A}']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100000,3'b000},// ['ALU{Y*A}']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100000,3'b000},// ['ALU{Y*A}']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100000,3'b000},// ['ALU{Y*A}']
	{2'b10,2'b00,6'b000000,5'b00011,2'b01,5'b11001,6'b100000,3'b000},// ['ALU{Y*A}', 'ALU{}->YA', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// D0 BNE
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// D1 TCALL 13
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101},// ['PCH->[SP]', 'SP//']
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100},// ['PCL->[SP]', 'SP//']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]->DR']
	{2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]:DR->PC']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// D2 CLR1 d.6
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010101,3'b000},// ['ALU{[AX]&~40}', 'ALU{}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// D3 BBC d.6
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// D4 MOV d+X, A
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+X->AL']
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b001},// ['A->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// D5 MOV !a+X, A
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b011000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'AL+X->AL', 'PC++']
	{2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AH+Carry->AH']
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b001},// ['A->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// D6 MOV !a+Y, A
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b011001,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'AL+X->AL', 'PC++']
	{2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AH+Carry->AH']
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b001},// ['A->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// D7 MOV {d}+Y, A
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR', 'AL+1->AL']
	{2'b00,2'b01,6'b011011,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->AH', 'DR+Y->AL']
	{2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AH+Carry->AH']
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b001},// ['A->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// D8 MOV d, X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00100,6'b000000,3'b001},// ['X->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// D9 MOV d+Y, X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b010001,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+Y->AL']
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00100,6'b000000,3'b001},// ['X->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// DA MOV d, YA
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]']
	{2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b001},// ['A->[AX]', 'AL+1->AL']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01000,6'b000000,3'b001},// ['Y->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// DB MOV d+X, Y
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+X->AL']
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01000,6'b000000,3'b001},// ['A->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// DC DEC Y
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00011,2'b11,5'b01001,6'b000010,3'b000},// ['ALU{Y-1}', 'ALU{}->Y', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// DD MOV A, Y
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00011,2'b01,5'b01001,6'b000000,3'b000},// ['ALU{Y}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// DE CBNE d+X, r
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+X->AL']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b010011,3'b000},// ['ALU{[AX]}']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// DF DAA
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00111,2'b01,5'b00000,6'b011110,3'b000},// ['ALU{A}->A', 'Flags']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// E0 CLRV
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b01000,2'b00,5'b00000,6'b000000,3'b000},// ['Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// E1 TCALL 14
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101},// ['PCH->[SP]', 'SP//']
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100},// ['PCL->[SP]', 'SP//']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]->DR']
	{2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]:DR->PC']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// E2 SET1 d.7
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010110,3'b000},// ['ALU{[AX]|80}', 'ALU{}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},	
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// E3 BBS d.7
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// E4 MOV A, d
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000000,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// E5 MOV A, !a
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'PC++']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000000,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// E6 MOV A, {X}
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100101,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['X->AL', 'P->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000000,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// E7 MOV A, {d+X}
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+X->AL']
	{2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR', 'AL+1->AL']
	{2'b00,2'b01,6'b011010,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->AH', 'DR->AL']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000000,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// E8 MOV A, #i
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00010,2'b01,5'b00000,6'b000000,3'b000},// ['ALU{[PC]}->A', 'PC++', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// E9 X, !a
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'PC++']
	{2'b10,2'b01,6'b000000,5'b00011,2'b10,5'b00000,6'b000000,3'b000},// ['ALU{[AX]}->X', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// EA NOT1 m.b
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]&1F->AH', '[PC]->DR', 'PC++']
	{2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b011011,3'b000},// ['ALU{[AX]}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// EB MOV Y, d
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b10,2'b01,6'b000000,5'b00011,2'b11,5'b00000,6'b000000,3'b000},// ['ALU{[AX]}->Y', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// EC Y, !a
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'PC++']
	{2'b10,2'b01,6'b000000,5'b00011,2'b11,5'b00000,6'b000000,3'b000},// ['ALU{[AX]}->Y', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// ED NOT C
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b01010,2'b00,5'b10100,6'b011100,3'b000},// ['C ^ 1']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// EE POP Y
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b10000,2'b00,5'b00000,6'b000000,3'b000},// ['SP++']
	{2'b00,2'b10,6'b000000,5'b00000,2'b11,5'b00000,6'b000000,3'b000},// ['[SP]->Y']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},//
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// EF SLEEP
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// F0 BEQ
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},	
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// F1 TCALL 15
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101},// ['PCH->[SP]', 'SP//']
	{2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100},// ['PCL->[SP]', 'SP//']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]->DR ']
	{2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000},// ['[VECT]:DR->PC ']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// F2 CLR1 d.7
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010101,3'b000},// ['ALU{[AX]&~80}', 'ALU{}->T']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// F3 BBC d.7
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// F4 MOV A, d+X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+X->AL']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000000,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// F5 MOV A, !a+X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b011000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'AL+X->AL', 'PC++']
	{2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AH+Carry->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000000,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// F6 MOV A, !a+Y
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'PC++']
	{2'b00,2'b00,6'b011001,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AH', 'AL+X->AL', 'PC++']
	{2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AH+Carry->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000000,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},	
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// F7 MOV A, {d}+Y
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->DR', 'AL+1->AL']
	{2'b00,2'b01,6'b011011,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->AH', 'DR+Y->AL']
	{2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AH+Carry->AH']
	{2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000000,3'b000},// ['ALU{[AX]}->A', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// F8 MOV X, d
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b10,2'b01,6'b000000,5'b00011,2'b10,5'b00000,6'b000000,3'b000},// ['ALU{[AX]}->X', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// F9 MOV X, d+Y
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b010001,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+Y->AL']
	{2'b10,2'b01,6'b000000,5'b00011,2'b10,5'b00000,6'b000000,3'b000},// ['ALU{[AX]}->X', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// FA MOV dd, ds
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b01,6'b000000,5'b00110,2'b00,5'b00000,6'b000000,3'b000},// ['[AX]->T']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001},// ['T->[AX]']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// FB MOV Y, d+X
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->AL', 'P->AH', 'PC++']
	{2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// ['AL+X->AL']
	{2'b10,2'b01,6'b000000,5'b00011,2'b11,5'b00000,6'b000000,3'b000},// ['ALU{[AX]}->Y', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// FC INC Y
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00011,2'b11,5'b01001,6'b000011,3'b000},// ['ALU{Y}->Y', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// FD MOV Y, A
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b10,2'b00,6'b000000,5'b00011,2'b11,5'b00001,6'b000000,3'b000},// ['ALU{A}->Y', 'Flags']
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// FE DBNZ Y, r
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b00,2'b00,6'b000000,5'b00000,2'b11,5'b01001,6'b000010,3'b000},// ['ALU{Y}->Y', 'Flags']
	{2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['[PC]->DR', 'PC++']
	{2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000},// ['PC+DR->PC']
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	// FF STOP
	{2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000},// ['PC++']
	{2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000},// []
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX},
	{2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX}    
} /* synthesis syn_ramstyle = "distributed_ram" */;

localparam ALUCtrl_r ALU_TAB[0:33] = '{
	{3'b110,4'b0011,1'b0,1'b0,1'b0},// 000000 LOAD
	{3'b100,4'b1011,1'b0,1'b1,1'b0},// 000001 DECW
	{3'b101,4'b1011,1'b0,1'b0,1'b0},// 000010 DEC 
	{3'b101,4'b1001,1'b0,1'b0,1'b0},// 000011 INC
	{3'b110,4'b0000,1'b0,1'b0,1'b0},// 000100 OR
	{3'b110,4'b0001,1'b0,1'b0,1'b0},// 000101 AND
	{3'b110,4'b0010,1'b0,1'b0,1'b0},// 000110 EOR
	{3'b110,4'b1000,1'b1,1'b0,1'b1},// 000111 ADC
	{3'b110,4'b1010,1'b1,1'b0,1'b1},// 001000 SBC
	{3'b100,4'b1001,1'b0,1'b1,1'b0},// 001001 INCW
	{3'b000,4'b0011,1'b0,1'b0,1'b1},// 001010 ASL
	{3'b010,4'b0011,1'b0,1'b0,1'b1},// 001011 LSR
	{3'b001,4'b0011,1'b0,1'b0,1'b1},// 001100 ROL
	{3'b011,4'b0011,1'b0,1'b0,1'b1},// 001101 ROR
	{3'b110,4'b0100,1'b0,1'b0,1'b0},// 001110 TCLR1
	{3'b110,4'b0101,1'b0,1'b0,1'b0},// 001111 TSET1
	{3'b110,4'b1011,1'b0,1'b1,1'b1},// 010000 CMPW
	{3'b110,4'b1001,1'b0,1'b0,1'b1},// 010001 ADD
	{3'b110,4'b1001,1'b1,1'b1,1'b1},// 010010 ADDW
	{3'b110,4'b1011,1'b0,1'b0,1'b1},// 010011 SUB/CMP
	{3'b110,4'b1011,1'b1,1'b1,1'b1},// 010100 SUBW
	{3'b111,4'b0001,1'b0,1'b0,1'b0},// 010101 CLR1
	{3'b110,4'b0000,1'b0,1'b0,1'b0},// 010110 SET1
	{3'b110,4'b0001,1'b0,1'b0,1'b0},// 010111 AND1
	{3'b111,4'b0001,1'b0,1'b0,1'b0},// 011000 NOT AND1
	{3'b110,4'b0000,1'b0,1'b0,1'b0},// 011001 OR1
	{3'b111,4'b0000,1'b0,1'b0,1'b0},// 011010 NOT OR1
	{3'b110,4'b0010,1'b0,1'b0,1'b0},// 011011 EOR1
	{3'b101,4'b0010,1'b0,1'b0,1'b0},// 011100 NOTC {C ^ 1}
	{3'b110,4'b0110,1'b0,1'b0,1'b0},// 011101 XCN
	{3'b110,4'b1100,1'b0,1'b0,1'b1},// 011110 DAA 
	{3'b110,4'b1101,1'b0,1'b0,1'b1},// 011111 DAS
	{3'b110,4'b1110,1'b0,1'b0,1'b0},// 100000 MUL 
	{3'b110,4'b1111,1'b1,1'b0,1'b0} // 100001 DIV
};

localparam RegCtrl_r REG_TAB[0:18] = '{
	{3'b000,2'b00,3'b000,2'b00},//00000
	{3'b001,2'b00,3'b000,2'b00},//00001 PC++
	{3'b001,2'b00,3'b001,2'b00},//00010 PC++, Flags
	{3'b000,2'b00,3'b001,2'b00},//00011 Flags
	{3'b000,2'b11,3'b000,2'b00},//00100 X->SP
	{3'b001,2'b00,3'b000,2'b01},//00101 [PC]->T, PC++
	{3'b000,2'b00,3'b000,2'b01},//00110 []->T
	{3'b000,2'b00,3'b001,2'b10},//00111 ALU{}->T, Flags
	{3'b000,2'b00,3'b100,2'b00},//01000 CLR/SET
	{3'b011,2'b00,3'b000,2'b00},//01001 PC+DR->PC
	{3'b000,2'b00,3'b101,2'b00},//01010 C change
	{3'b000,2'b00,3'b000,2'b10},//01011 ALU{}->T
	{3'b010,2'b00,3'b000,2'b00},//01100 []:DR->PC
	{3'b000,2'b10,3'b000,2'b00},//01101 Reg->[SP], SP//
	{3'b100,2'b00,3'b000,2'b00},//01110 AX->PC
	{3'b000,2'b00,3'b010,2'b00},//01111 1->B
	{3'b000,2'b01,3'b000,2'b00},//10000 SP++
	{3'b000,2'b00,3'b011,2'b00},//10001 []->PSW
	{3'b101,2'b00,3'b000,2'b00} //10010 FF:AL->PC
};

MicroInst_r MI;
ALUCtrl_r ALUFlags;
RegCtrl_r R;

assign ALUFlags = ALU_TAB[MI.ALUCtrl];
assign R = REG_TAB[MI.regMode];

always @(posedge CLK) begin
    if (~RST_N)
        MI <= {2'b0, 2'b0, 6'b0, 5'b1, 2'b0, 5'b0, 6'b0, 3'b0};
    else 
        if (EN)
            MI <= M_TAB[{IR, STATE}];
end

assign M = {ALUFlags, 
            MI.stateCtrl, 
            MI.addrBus, 
            MI.addrCtrl,
            R.loadPC,
            R.loadSP, 
            MI.regAXY, 
            R.loadP, 
            R.loadT,
            MI.busCtrl,
            MI.outBus};

endmodule